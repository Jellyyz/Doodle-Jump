module LFSR(
    input 
    input 
    output
); 


endmodule 


module sixteen_bit_register(
    input Clk; 
    input D; 
    output Q; 
); 


endmodule 